// Automatically generated Verilog-2005
module HeapSort_testInput_14(// clock
                            system1000
                            ,// asynchronous reset: active low
                            system1000_rstn
                            ,topLet_o);
  input system1000;
  input system1000_rstn;
  output [160:0] topLet_o;
  HeapSort_stimuliGeneratorzm_15 HeapSort_stimuliGeneratorzm_15_topLet_o
  (.bodyVar_o (topLet_o)
  ,.system1000 (system1000)
  ,.system1000_rstn (system1000_rstn));
endmodule
