-- Automatically generated VHDL-2002
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;
use std.textio.all;
use work.all;
use work.Path_types.all;

entity Path_testInput_15 is
  port(topLet_o : out std_logic_vector(64 downto 0));
end;

architecture structural of Path_testInput_15 is
begin
  topLet_o <= std_logic_vector'("1" & (std_logic_vector(unsigned'("0000000000000100"))
                                       & std_logic_vector(unsigned'("0000000000000100"))
                                       & std_logic_vector(unsigned'("0000000000000011"))
                                       & std_logic_vector(unsigned'("0000000000001111"))));
end;
