// Automatically generated Verilog-2005
module Path_testInput_15(topLet_o);
  output [64:0] topLet_o;
  assign topLet_o = {1'b1,{16'd4
                          ,16'd4
                          ,16'd3
                          ,16'd15}};
endmodule
